--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   18:39:11 04/30/2020
-- Design Name:   
-- Module Name:   /home/janfrolka/projekt/druhytestbench7SEG.vhd
-- Project Name:  projekt
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: hex_to_7seg
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY druhytestbench7SEG IS
END druhytestbench7SEG;
 
ARCHITECTURE behavior OF druhytestbench7SEG IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT hex_to_7seg
    PORT(
         hex_i : IN  std_logic_vector(3 downto 0);
         seg_o : OUT  std_logic_vector(6 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal hex_i : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal seg_o : std_logic_vector(6 downto 0);
   -- No clocks detected in port list. Replace <clock> below with 
   -- appropriate port name 
 
   --constant clock_period : time := 100 ms;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: hex_to_7seg PORT MAP (
          hex_i => hex_i,
          seg_o => seg_o
        );

   -- Clock process definitions
--   clock_process :process
--   begin
--		clock <= '0';
--		wait for clock_period/2;
--		clock <= '1';
--		wait for clock_period/2;
--   end process;
 

   -- Stimulus process
   stim_proc: process
   begin		
      -- hold reset state for 100 ns.
      wait for 100 ns;	

      --wait for clock_period*10;

      -- insert stimulus here 
		hex_i <= "1001";

      wait;
   end process;

END;
